module tb;
`include "readme.txt"

endmodule